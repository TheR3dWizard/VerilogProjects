module speed (input clk,rst,input [7:0] force)