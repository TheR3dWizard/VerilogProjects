module comparison